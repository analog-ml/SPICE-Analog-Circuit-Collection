Tan_CLIA_Pin_3


*-----------------------------------------------------------
* Model LIB definition
*-----------------------------------------------------------
.param mc_mm_switch=0
.param mc_pr_switch=0
*.include /home/pham/shared_files/sky130_pdk/libs.tech/ngspice/corners/tt.spice
*.include /home/pham/shared_files/sky130_pdk/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
*.include /home/pham/shared_files/sky130_pdk/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
*.include /home/pham/shared_files/sky130_pdk/libs.tech/ngspice/corners/tt/specialized_cells.spice
.lib /home/pham/shared_files/sky130_pdk/libs.tech/ngspice/sky130.lib.spice tt

* Fixed PARAM
*-----------------------------------------------------------
.PARAM supply_voltage = 1.8
.PARAM VCM_ratio = 0.4


* Tunable PARAM
*-----------------------------------------------------------
.PARAM
+ MOSFET_5_2_L_LOAD1_PMOS=1 MOSFET_5_2_M_LOAD1_PMOS=117 
+ MOSFET_5_2_W_LOAD1_PMOS=1 CURRENT_0_BIAS=630n 
+ MOSFET_0_8_L_BIASCM_PMOS=1 MOSFET_0_8_M_BIASCM_PMOS=200 
+ MOSFET_0_8_W_BIASCM_PMOS=1 MOSFET_17_7_L_BIASCM_NMOS=1 
+ MOSFET_17_7_M_BIASCM_NMOS=1 MOSFET_17_7_W_BIASCM_NMOS=0.500 
+ MOSFET_68_1_L_gmf_PMOS=0.500 MOSFET_68_1_M_gmf_PMOS=6 
+ MOSFET_68_1_W_gmf_PMOS=1 MOSFET_69_1_L_gm3_NMOS=0.900 
+ MOSFET_69_1_M_gm3_NMOS=3 MOSFET_69_1_W_gm3_NMOS=1 
+ MOSFET_70_1_L_gm21_PMOS=0.480 MOSFET_70_1_M_gm21_PMOS=2 
+ MOSFET_70_1_W_gm21_PMOS=1 MOSFET_71_1_L_gm23_NMOS=1 
+ MOSFET_71_1_M_gm23_NMOS=1 MOSFET_71_1_W_gm23_NMOS=0.453 
+ MOSFET_8_2_L_gm1_PMOS=1 MOSFET_8_2_M_gm1_PMOS=100 
+ MOSFET_8_2_W_gm1_PMOS=1 RESISTOR_0=247.56K CAPACITOR_0=347f 
+ CAPACITOR_1=240f CLOAD=560p VCM=300m 


.subckt tan_clia_pin_3 GNDA VDDA VINN VINP VOUT
xm73 net5 DM_1 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_0_8_L_BIASCM_PMOS' w='MOSFET_0_8_W_BIASCM_PMOS*1' m='12*MOSFET_0_8_M_BIASCM_PMOS'
xm70 net3 net050 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_70_1_L_gm21_PMOS' w='MOSFET_70_1_W_gm21_PMOS*1' m='MOSFET_70_1_M_gm21_PMOS'
xm2 DM_1 DM_1 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_0_8_L_BIASCM_PMOS' w='MOSFET_0_8_W_BIASCM_PMOS*1' m='MOSFET_0_8_M_BIASCM_PMOS*4'
xm68 VOUT net050 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_68_1_L_gmf_PMOS' w='MOSFET_68_1_W_gmf_PMOS*1' m='MOSFET_68_1_M_gmf_PMOS'
xm6 net050 VOUTN VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_5_2_L_LOAD1_PMOS' w='MOSFET_5_2_W_LOAD1_PMOS*1' m='MOSFET_5_2_M_LOAD1_PMOS'
xm5 VOUTN VOUTN VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_5_2_L_LOAD1_PMOS' w='MOSFET_5_2_W_LOAD1_PMOS*1' m='MOSFET_5_2_M_LOAD1_PMOS'
xm9 net8 VINP net31 net31 sky130_fd_pr__pfet_01v8 l='MOSFET_8_2_L_gm1_PMOS' w='MOSFET_8_2_W_gm1_PMOS*1' m='MOSFET_8_2_M_gm1_PMOS'
xm8 DM_2 VINN net31 net31 sky130_fd_pr__pfet_01v8 l='MOSFET_8_2_L_gm1_PMOS' w='MOSFET_8_2_W_gm1_PMOS*1' m='MOSFET_8_2_M_gm1_PMOS'
xm4 net31 net1 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_0_8_L_BIASCM_PMOS' w='MOSFET_0_8_W_BIASCM_PMOS*1' m='8*MOSFET_0_8_M_BIASCM_PMOS'
xm3 VB3 net1 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_0_8_L_BIASCM_PMOS' w='MOSFET_0_8_W_BIASCM_PMOS*1' m='MOSFET_0_8_M_BIASCM_PMOS*4'
xm1 VB4 net1 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_0_8_L_BIASCM_PMOS' w='MOSFET_0_8_W_BIASCM_PMOS*1' m='MOSFET_0_8_M_BIASCM_PMOS*4'
xm0 net1 net1 VDDA VDDA sky130_fd_pr__pfet_01v8 l='MOSFET_0_8_L_BIASCM_PMOS' w='MOSFET_0_8_W_BIASCM_PMOS*1' m='MOSFET_0_8_M_BIASCM_PMOS*4'
xm72 net5 net3 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_71_1_L_gm23_NMOS' w='MOSFET_71_1_W_gm23_NMOS*1' m='MOSFET_71_1_M_gm23_NMOS*3'
xm61 net3 VB4 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*6'
xm71 net3 net3 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_71_1_L_gm23_NMOS' w='MOSFET_71_1_W_gm23_NMOS*1' m='MOSFET_71_1_M_gm23_NMOS'
xm19 DM_2 VB4 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*12'
xm15 VOUTN VB3 DM_2 GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*8'
xm20 net8 VB4 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*12'
xm16 net050 VB3 net8 GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*8'
xm18 net7 VB4 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*4'
xm12 VB4 VB3 net6 GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*4'
xm13 DM_1 VB3 net7 GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*4'
xm17 net6 VB4 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS*4'
xm69 VOUT net5 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_69_1_L_gm3_NMOS' w='MOSFET_69_1_W_gm3_NMOS*1' m='MOSFET_69_1_M_gm3_NMOS'
xm14 VB3 VB3 GNDA GNDA sky130_fd_pr__nfet_01v8 l='MOSFET_17_7_L_BIASCM_NMOS' w='MOSFET_17_7_W_BIASCM_NMOS*1' m='MOSFET_17_7_M_BIASCM_NMOS'
I0 net1 GNDA 'CURRENT_0_BIAS'
C1 net8 VOUT 'CAPACITOR_1'
C0 net2 GNDA 'CAPACITOR_0'
R0 net5 net2 'RESISTOR_0'
.ends tan_clia_pin_3

*-----------------------------------------------------------
* Parameter definition
*-----------------------------------------------------------




V1 vdd 0 'supply_voltage'
V2 vss 0 0 

Vindc opin 0 'supply_voltage*VCM_ratio'
Vin signal_in 0 dc 'supply_voltage*VCM_ratio' ac 1 sin('supply_voltage*VCM_ratio' 100m 500)

Lfb opout opout_dc 1T
Cin opout_dc signal_in 1T

x1 vss vdd opout_dc opin opout  tan_clia_pin_3
Cload1 opout 0 'CLOAD'


.ac dec 10 1 10G

.control
    run
    set units=degrees
    set wr_vecnames
    option numdgt=7
    
    meas ac gain_bandwidth_product when vdb(opout)=0
    meas ac phase_margin find vp(opout) when vdb(opout)=0
    wrdata CLIA_GBW_PM  gain_bandwidth_product phase_margin 

    wrdata ac.csv v(opout)
    op
    wrdata dc.csv i(V1)

    set filetype=ascii
.endc

.end