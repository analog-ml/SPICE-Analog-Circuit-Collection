let gmbs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[gm]
let gds_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[vth]
let id_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[id]
let ibd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[igs]
let igd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[igd]
let igb_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cds]
let csg_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[csg]
let csd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[csd]
let css_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[css]
let cgb_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM11=@m.x1.xm11.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[gm]
let gds_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[vth]
let id_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[id]
let ibd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[igs]
let igd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[igd]
let igb_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cds]
let csg_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[csg]
let csd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[csd]
let css_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[css]
let cgb_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM7=@m.x1.xm7.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[gm]
let gds_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[vth]
let id_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[id]
let ibd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[igs]
let igd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[igd]
let igb_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cds]
let csg_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[csg]
let csd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[csd]
let css_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[css]
let cgb_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM10=@m.x1.xm10.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[gm]
let gds_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[vth]
let id_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[id]
let ibd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[igs]
let igd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[igd]
let igb_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cds]
let csg_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[csg]
let csd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[csd]
let css_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[css]
let cgb_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM6=@m.x1.xm6.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[gm]
let gds_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[vth]
let id_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[id]
let ibd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[igs]
let igd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[igd]
let igb_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cds]
let csg_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[csg]
let csd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[csd]
let css_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[css]
let cgb_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM5=@m.x1.xm5.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[gm]
let gds_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[vth]
let id_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[id]
let ibd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[igs]
let igd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[igd]
let igb_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cds]
let csg_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[csg]
let csd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[csd]
let css_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[css]
let cgb_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM9=@m.x1.xm9.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[gm]
let gds_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[vth]
let id_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[id]
let ibd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[igs]
let igd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[igd]
let igb_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cds]
let csg_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[csg]
let csd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[csd]
let css_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[css]
let cgb_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM8=@m.x1.xm8.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[gm]
let gds_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[vth]
let id_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[id]
let ibd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[igs]
let igd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[igd]
let igb_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cds]
let csg_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[csg]
let csd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[csd]
let css_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[css]
let cgb_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM4=@m.x1.xm4.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[gm]
let gds_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[vth]
let id_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[id]
let ibd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[igs]
let igd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[igd]
let igb_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cds]
let csg_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[csg]
let csd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[csd]
let css_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[css]
let cgb_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM3=@m.x1.xm3.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[gm]
let gds_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[vth]
let id_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[id]
let ibd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[igs]
let igd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[igd]
let igb_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cds]
let csg_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[csg]
let csd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[csd]
let css_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[css]
let cgb_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM2=@m.x1.xm2.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[gm]
let gds_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[vth]
let id_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[id]
let ibd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[igs]
let igd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[igd]
let igb_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cds]
let csg_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[csg]
let csd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[csd]
let css_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[css]
let cgb_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM1=@m.x1.xm1.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[gmbs]
let gm_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[gm]
let gds_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[gds]
let vdsat_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[vdsat]
let vth_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[vth]
let id_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[id]
let ibd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[ibd]
let ibs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[ibs]
let gbd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[gbd]
let gbs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[gbs]
let isub_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[isub]
let igidl_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[igidl]
let igisl_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[igisl]
let igs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[igs]
let igd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[igd]
let igb_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[igb]
let igcs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[igcs]
let vbs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[vbs]
let vgs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[vgs]
let vds_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[vds]
let cgg_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cgg]
let cgs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cgs]
let cgd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cgd]
let cbg_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cbg]
let cbd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cbd]
let cbs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cbs]
let cdg_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cdg]
let cdd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cdd]
let cds_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cds]
let csg_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[csg]
let csd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[csd]
let css_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[css]
let cgb_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cgb]
let cdb_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cdb]
let csb_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[csb]
let cbb_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[cbb]
let capbd_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[capbd]
let capbs_XM0=@m.x1.xm0.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[gm]
let gds_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[vth]
let id_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[id]
let ibd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[igs]
let igd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[igd]
let igb_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cds]
let csg_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[csg]
let csd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[csd]
let css_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[css]
let cgb_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM23=@m.x1.xm23.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[gm]
let gds_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[vth]
let id_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[id]
let ibd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[igs]
let igd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[igd]
let igb_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cds]
let csg_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[csg]
let csd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[csd]
let css_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[css]
let cgb_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM22=@m.x1.xm22.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[gm]
let gds_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[vth]
let id_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[id]
let ibd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[igs]
let igd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[igd]
let igb_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cds]
let csg_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[csg]
let csd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[csd]
let css_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[css]
let cgb_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM21=@m.x1.xm21.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[gm]
let gds_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[vth]
let id_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[id]
let ibd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[igs]
let igd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[igd]
let igb_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cds]
let csg_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[csg]
let csd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[csd]
let css_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[css]
let cgb_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM19=@m.x1.xm19.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[gm]
let gds_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[vth]
let id_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[id]
let ibd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[igs]
let igd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[igd]
let igb_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cds]
let csg_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[csg]
let csd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[csd]
let css_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[css]
let cgb_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM15=@m.x1.xm15.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[gm]
let gds_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[vth]
let id_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[id]
let ibd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[igs]
let igd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[igd]
let igb_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cds]
let csg_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[csg]
let csd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[csd]
let css_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[css]
let cgb_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM20=@m.x1.xm20.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[gm]
let gds_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[vth]
let id_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[id]
let ibd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[igs]
let igd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[igd]
let igb_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cds]
let csg_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[csg]
let csd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[csd]
let css_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[css]
let cgb_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM16=@m.x1.xm16.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[gm]
let gds_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[vth]
let id_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[id]
let ibd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[igs]
let igd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[igd]
let igb_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cds]
let csg_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[csg]
let csd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[csd]
let css_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[css]
let cgb_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM17=@m.x1.xm17.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[gm]
let gds_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[vth]
let id_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[id]
let ibd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[igs]
let igd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[igd]
let igb_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cds]
let csg_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[csg]
let csd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[csd]
let css_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[css]
let cgb_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM14=@m.x1.xm14.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[gm]
let gds_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[vth]
let id_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[id]
let ibd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[igs]
let igd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[igd]
let igb_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cds]
let csg_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[csg]
let csd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[csd]
let css_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[css]
let cgb_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM12=@m.x1.xm12.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[gm]
let gds_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[vth]
let id_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[id]
let ibd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[igs]
let igd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[igd]
let igb_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cds]
let csg_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[csg]
let csd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[csd]
let css_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[css]
let cgb_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM18=@m.x1.xm18.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[gmbs]
let gm_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[gm]
let gds_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[gds]
let vdsat_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[vdsat]
let vth_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[vth]
let id_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[id]
let ibd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[ibd]
let ibs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[ibs]
let gbd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[gbd]
let gbs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[gbs]
let isub_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[isub]
let igidl_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[igidl]
let igisl_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[igisl]
let igs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[igs]
let igd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[igd]
let igb_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[igb]
let igcs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[igcs]
let vbs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[vbs]
let vgs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[vgs]
let vds_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[vds]
let cgg_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cgg]
let cgs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cgs]
let cgd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cgd]
let cbg_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cbg]
let cbd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cbd]
let cbs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cbs]
let cdg_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cdg]
let cdd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cdd]
let cds_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cds]
let csg_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[csg]
let csd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[csd]
let css_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[css]
let cgb_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cgb]
let cdb_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cdb]
let csb_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[csb]
let cbb_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[cbb]
let capbd_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[capbd]
let capbs_XM13=@m.x1.xm13.msky130_fd_pr__nfet_01v8[capbs]

let capacitance_XC0=@c.x1.xc0.c1[capacitance]
let cap_XC0=@c.x1.xc0.c1[cap]
let c_XC0=@c.x1.xc0.c1[c]
let ic_XC0=@c.x1.xc0.c1[ic]
let temp_XC0=@c.x1.xc0.c1[temp]
let dtemp_XC0=@c.x1.xc0.c1[dtemp]
let w_XC0=@c.x1.xc0.c1[w]
let l_XC0=@c.x1.xc0.c1[l]
let m_XC0=@c.x1.xc0.c1[m]
let scale_XC0=@c.x1.xc0.c1[scale]
let i_XC0=@c.x1.xc0.c1[i]
let p_XC0=@c.x1.xc0.c1[p]
let sens_dc_XC0=@c.x1.xc0.c1[sens_dc]
let sens_real_XC0=@c.x1.xc0.c1[sens_real]
let sens_imag_XC0=@c.x1.xc0.c1[sens_imag]
let sens_mag_XC0=@c.x1.xc0.c1[sens_mag]
let sens_ph_XC0=@c.x1.xc0.c1[sens_ph]
let sens_cplx_XC0=@c.x1.xc0.c1[sens_cplx]

let capacitance_XC1=@c.x1.xc1.c1[capacitance]
let cap_XC1=@c.x1.xc1.c1[cap]
let c_XC1=@c.x1.xc1.c1[c]
let ic_XC1=@c.x1.xc1.c1[ic]
let temp_XC1=@c.x1.xc1.c1[temp]
let dtemp_XC1=@c.x1.xc1.c1[dtemp]
let w_XC1=@c.x1.xc1.c1[w]
let l_XC1=@c.x1.xc1.c1[l]
let m_XC1=@c.x1.xc1.c1[m]
let scale_XC1=@c.x1.xc1.c1[scale]
let i_XC1=@c.x1.xc1.c1[i]
let p_XC1=@c.x1.xc1.c1[p]
let sens_dc_XC1=@c.x1.xc1.c1[sens_dc]
let sens_real_XC1=@c.x1.xc1.c1[sens_real]
let sens_imag_XC1=@c.x1.xc1.c1[sens_imag]
let sens_mag_XC1=@c.x1.xc1.c1[sens_mag]
let sens_ph_XC1=@c.x1.xc1.c1[sens_ph]
let sens_cplx_XC1=@c.x1.xc1.c1[sens_cplx]

write Leung_NMCF_region gmbs_XM11 gm_XM11 gds_XM11 vdsat_XM11 vth_XM11 id_XM11 ibd_XM11 ibs_XM11 gbd_XM11 gbs_XM11 isub_XM11 igidl_XM11 igisl_XM11 igs_XM11 igd_XM11 igb_XM11 igcs_XM11 vbs_XM11 vgs_XM11 vds_XM11 cgg_XM11 cgs_XM11 cgd_XM11 cbg_XM11 cbd_XM11 cbs_XM11 cdg_XM11 cdd_XM11 cds_XM11 csg_XM11 csd_XM11 css_XM11 cgb_XM11 cdb_XM11 csb_XM11 cbb_XM11 capbd_XM11 capbs_XM11 gmbs_XM7 gm_XM7 gds_XM7 vdsat_XM7 vth_XM7 id_XM7 ibd_XM7 ibs_XM7 gbd_XM7 gbs_XM7 isub_XM7 igidl_XM7 igisl_XM7 igs_XM7 igd_XM7 igb_XM7 igcs_XM7 vbs_XM7 vgs_XM7 vds_XM7 cgg_XM7 cgs_XM7 cgd_XM7 cbg_XM7 cbd_XM7 cbs_XM7 cdg_XM7 cdd_XM7 cds_XM7 csg_XM7 csd_XM7 css_XM7 cgb_XM7 cdb_XM7 csb_XM7 cbb_XM7 capbd_XM7 capbs_XM7 gmbs_XM10 gm_XM10 gds_XM10 vdsat_XM10 vth_XM10 id_XM10 ibd_XM10 ibs_XM10 gbd_XM10 gbs_XM10 isub_XM10 igidl_XM10 igisl_XM10 igs_XM10 igd_XM10 igb_XM10 igcs_XM10 vbs_XM10 vgs_XM10 vds_XM10 cgg_XM10 cgs_XM10 cgd_XM10 cbg_XM10 cbd_XM10 cbs_XM10 cdg_XM10 cdd_XM10 cds_XM10 csg_XM10 csd_XM10 css_XM10 cgb_XM10 cdb_XM10 csb_XM10 cbb_XM10 capbd_XM10 capbs_XM10 gmbs_XM6 gm_XM6 gds_XM6 vdsat_XM6 vth_XM6 id_XM6 ibd_XM6 ibs_XM6 gbd_XM6 gbs_XM6 isub_XM6 igidl_XM6 igisl_XM6 igs_XM6 igd_XM6 igb_XM6 igcs_XM6 vbs_XM6 vgs_XM6 vds_XM6 cgg_XM6 cgs_XM6 cgd_XM6 cbg_XM6 cbd_XM6 cbs_XM6 cdg_XM6 cdd_XM6 cds_XM6 csg_XM6 csd_XM6 css_XM6 cgb_XM6 cdb_XM6 csb_XM6 cbb_XM6 capbd_XM6 capbs_XM6 gmbs_XM5 gm_XM5 gds_XM5 vdsat_XM5 vth_XM5 id_XM5 ibd_XM5 ibs_XM5 gbd_XM5 gbs_XM5 isub_XM5 igidl_XM5 igisl_XM5 igs_XM5 igd_XM5 igb_XM5 igcs_XM5 vbs_XM5 vgs_XM5 vds_XM5 cgg_XM5 cgs_XM5 cgd_XM5 cbg_XM5 cbd_XM5 cbs_XM5 cdg_XM5 cdd_XM5 cds_XM5 csg_XM5 csd_XM5 css_XM5 cgb_XM5 cdb_XM5 csb_XM5 cbb_XM5 capbd_XM5 capbs_XM5 gmbs_XM9 gm_XM9 gds_XM9 vdsat_XM9 vth_XM9 id_XM9 ibd_XM9 ibs_XM9 gbd_XM9 gbs_XM9 isub_XM9 igidl_XM9 igisl_XM9 igs_XM9 igd_XM9 igb_XM9 igcs_XM9 vbs_XM9 vgs_XM9 vds_XM9 cgg_XM9 cgs_XM9 cgd_XM9 cbg_XM9 cbd_XM9 cbs_XM9 cdg_XM9 cdd_XM9 cds_XM9 csg_XM9 csd_XM9 css_XM9 cgb_XM9 cdb_XM9 csb_XM9 cbb_XM9 capbd_XM9 capbs_XM9 gmbs_XM8 gm_XM8 gds_XM8 vdsat_XM8 vth_XM8 id_XM8 ibd_XM8 ibs_XM8 gbd_XM8 gbs_XM8 isub_XM8 igidl_XM8 igisl_XM8 igs_XM8 igd_XM8 igb_XM8 igcs_XM8 vbs_XM8 vgs_XM8 vds_XM8 cgg_XM8 cgs_XM8 cgd_XM8 cbg_XM8 cbd_XM8 cbs_XM8 cdg_XM8 cdd_XM8 cds_XM8 csg_XM8 csd_XM8 css_XM8 cgb_XM8 cdb_XM8 csb_XM8 cbb_XM8 capbd_XM8 capbs_XM8 gmbs_XM4 gm_XM4 gds_XM4 vdsat_XM4 vth_XM4 id_XM4 ibd_XM4 ibs_XM4 gbd_XM4 gbs_XM4 isub_XM4 igidl_XM4 igisl_XM4 igs_XM4 igd_XM4 igb_XM4 igcs_XM4 vbs_XM4 vgs_XM4 vds_XM4 cgg_XM4 cgs_XM4 cgd_XM4 cbg_XM4 cbd_XM4 cbs_XM4 cdg_XM4 cdd_XM4 cds_XM4 csg_XM4 csd_XM4 css_XM4 cgb_XM4 cdb_XM4 csb_XM4 cbb_XM4 capbd_XM4 capbs_XM4 gmbs_XM3 gm_XM3 gds_XM3 vdsat_XM3 vth_XM3 id_XM3 ibd_XM3 ibs_XM3 gbd_XM3 gbs_XM3 isub_XM3 igidl_XM3 igisl_XM3 igs_XM3 igd_XM3 igb_XM3 igcs_XM3 vbs_XM3 vgs_XM3 vds_XM3 cgg_XM3 cgs_XM3 cgd_XM3 cbg_XM3 cbd_XM3 cbs_XM3 cdg_XM3 cdd_XM3 cds_XM3 csg_XM3 csd_XM3 css_XM3 cgb_XM3 cdb_XM3 csb_XM3 cbb_XM3 capbd_XM3 capbs_XM3 gmbs_XM2 gm_XM2 gds_XM2 vdsat_XM2 vth_XM2 id_XM2 ibd_XM2 ibs_XM2 gbd_XM2 gbs_XM2 isub_XM2 igidl_XM2 igisl_XM2 igs_XM2 igd_XM2 igb_XM2 igcs_XM2 vbs_XM2 vgs_XM2 vds_XM2 cgg_XM2 cgs_XM2 cgd_XM2 cbg_XM2 cbd_XM2 cbs_XM2 cdg_XM2 cdd_XM2 cds_XM2 csg_XM2 csd_XM2 css_XM2 cgb_XM2 cdb_XM2 csb_XM2 cbb_XM2 capbd_XM2 capbs_XM2 gmbs_XM1 gm_XM1 gds_XM1 vdsat_XM1 vth_XM1 id_XM1 ibd_XM1 ibs_XM1 gbd_XM1 gbs_XM1 isub_XM1 igidl_XM1 igisl_XM1 igs_XM1 igd_XM1 igb_XM1 igcs_XM1 vbs_XM1 vgs_XM1 vds_XM1 cgg_XM1 cgs_XM1 cgd_XM1 cbg_XM1 cbd_XM1 cbs_XM1 cdg_XM1 cdd_XM1 cds_XM1 csg_XM1 csd_XM1 css_XM1 cgb_XM1 cdb_XM1 csb_XM1 cbb_XM1 capbd_XM1 capbs_XM1 gmbs_XM0 gm_XM0 gds_XM0 vdsat_XM0 vth_XM0 id_XM0 ibd_XM0 ibs_XM0 gbd_XM0 gbs_XM0 isub_XM0 igidl_XM0 igisl_XM0 igs_XM0 igd_XM0 igb_XM0 igcs_XM0 vbs_XM0 vgs_XM0 vds_XM0 cgg_XM0 cgs_XM0 cgd_XM0 cbg_XM0 cbd_XM0 cbs_XM0 cdg_XM0 cdd_XM0 cds_XM0 csg_XM0 csd_XM0 css_XM0 cgb_XM0 cdb_XM0 csb_XM0 cbb_XM0 capbd_XM0 capbs_XM0 gmbs_XM23 gm_XM23 gds_XM23 vdsat_XM23 vth_XM23 id_XM23 ibd_XM23 ibs_XM23 gbd_XM23 gbs_XM23 isub_XM23 igidl_XM23 igisl_XM23 igs_XM23 igd_XM23 igb_XM23 igcs_XM23 vbs_XM23 vgs_XM23 vds_XM23 cgg_XM23 cgs_XM23 cgd_XM23 cbg_XM23 cbd_XM23 cbs_XM23 cdg_XM23 cdd_XM23 cds_XM23 csg_XM23 csd_XM23 css_XM23 cgb_XM23 cdb_XM23 csb_XM23 cbb_XM23 capbd_XM23 capbs_XM23 gmbs_XM22 gm_XM22 gds_XM22 vdsat_XM22 vth_XM22 id_XM22 ibd_XM22 ibs_XM22 gbd_XM22 gbs_XM22 isub_XM22 igidl_XM22 igisl_XM22 igs_XM22 igd_XM22 igb_XM22 igcs_XM22 vbs_XM22 vgs_XM22 vds_XM22 cgg_XM22 cgs_XM22 cgd_XM22 cbg_XM22 cbd_XM22 cbs_XM22 cdg_XM22 cdd_XM22 cds_XM22 csg_XM22 csd_XM22 css_XM22 cgb_XM22 cdb_XM22 csb_XM22 cbb_XM22 capbd_XM22 capbs_XM22 gmbs_XM21 gm_XM21 gds_XM21 vdsat_XM21 vth_XM21 id_XM21 ibd_XM21 ibs_XM21 gbd_XM21 gbs_XM21 isub_XM21 igidl_XM21 igisl_XM21 igs_XM21 igd_XM21 igb_XM21 igcs_XM21 vbs_XM21 vgs_XM21 vds_XM21 cgg_XM21 cgs_XM21 cgd_XM21 cbg_XM21 cbd_XM21 cbs_XM21 cdg_XM21 cdd_XM21 cds_XM21 csg_XM21 csd_XM21 css_XM21 cgb_XM21 cdb_XM21 csb_XM21 cbb_XM21 capbd_XM21 capbs_XM21 gmbs_XM19 gm_XM19 gds_XM19 vdsat_XM19 vth_XM19 id_XM19 ibd_XM19 ibs_XM19 gbd_XM19 gbs_XM19 isub_XM19 igidl_XM19 igisl_XM19 igs_XM19 igd_XM19 igb_XM19 igcs_XM19 vbs_XM19 vgs_XM19 vds_XM19 cgg_XM19 cgs_XM19 cgd_XM19 cbg_XM19 cbd_XM19 cbs_XM19 cdg_XM19 cdd_XM19 cds_XM19 csg_XM19 csd_XM19 css_XM19 cgb_XM19 cdb_XM19 csb_XM19 cbb_XM19 capbd_XM19 capbs_XM19 gmbs_XM15 gm_XM15 gds_XM15 vdsat_XM15 vth_XM15 id_XM15 ibd_XM15 ibs_XM15 gbd_XM15 gbs_XM15 isub_XM15 igidl_XM15 igisl_XM15 igs_XM15 igd_XM15 igb_XM15 igcs_XM15 vbs_XM15 vgs_XM15 vds_XM15 cgg_XM15 cgs_XM15 cgd_XM15 cbg_XM15 cbd_XM15 cbs_XM15 cdg_XM15 cdd_XM15 cds_XM15 csg_XM15 csd_XM15 css_XM15 cgb_XM15 cdb_XM15 csb_XM15 cbb_XM15 capbd_XM15 capbs_XM15 gmbs_XM20 gm_XM20 gds_XM20 vdsat_XM20 vth_XM20 id_XM20 ibd_XM20 ibs_XM20 gbd_XM20 gbs_XM20 isub_XM20 igidl_XM20 igisl_XM20 igs_XM20 igd_XM20 igb_XM20 igcs_XM20 vbs_XM20 vgs_XM20 vds_XM20 cgg_XM20 cgs_XM20 cgd_XM20 cbg_XM20 cbd_XM20 cbs_XM20 cdg_XM20 cdd_XM20 cds_XM20 csg_XM20 csd_XM20 css_XM20 cgb_XM20 cdb_XM20 csb_XM20 cbb_XM20 capbd_XM20 capbs_XM20 gmbs_XM16 gm_XM16 gds_XM16 vdsat_XM16 vth_XM16 id_XM16 ibd_XM16 ibs_XM16 gbd_XM16 gbs_XM16 isub_XM16 igidl_XM16 igisl_XM16 igs_XM16 igd_XM16 igb_XM16 igcs_XM16 vbs_XM16 vgs_XM16 vds_XM16 cgg_XM16 cgs_XM16 cgd_XM16 cbg_XM16 cbd_XM16 cbs_XM16 cdg_XM16 cdd_XM16 cds_XM16 csg_XM16 csd_XM16 css_XM16 cgb_XM16 cdb_XM16 csb_XM16 cbb_XM16 capbd_XM16 capbs_XM16 gmbs_XM17 gm_XM17 gds_XM17 vdsat_XM17 vth_XM17 id_XM17 ibd_XM17 ibs_XM17 gbd_XM17 gbs_XM17 isub_XM17 igidl_XM17 igisl_XM17 igs_XM17 igd_XM17 igb_XM17 igcs_XM17 vbs_XM17 vgs_XM17 vds_XM17 cgg_XM17 cgs_XM17 cgd_XM17 cbg_XM17 cbd_XM17 cbs_XM17 cdg_XM17 cdd_XM17 cds_XM17 csg_XM17 csd_XM17 css_XM17 cgb_XM17 cdb_XM17 csb_XM17 cbb_XM17 capbd_XM17 capbs_XM17 gmbs_XM14 gm_XM14 gds_XM14 vdsat_XM14 vth_XM14 id_XM14 ibd_XM14 ibs_XM14 gbd_XM14 gbs_XM14 isub_XM14 igidl_XM14 igisl_XM14 igs_XM14 igd_XM14 igb_XM14 igcs_XM14 vbs_XM14 vgs_XM14 vds_XM14 cgg_XM14 cgs_XM14 cgd_XM14 cbg_XM14 cbd_XM14 cbs_XM14 cdg_XM14 cdd_XM14 cds_XM14 csg_XM14 csd_XM14 css_XM14 cgb_XM14 cdb_XM14 csb_XM14 cbb_XM14 capbd_XM14 capbs_XM14 gmbs_XM12 gm_XM12 gds_XM12 vdsat_XM12 vth_XM12 id_XM12 ibd_XM12 ibs_XM12 gbd_XM12 gbs_XM12 isub_XM12 igidl_XM12 igisl_XM12 igs_XM12 igd_XM12 igb_XM12 igcs_XM12 vbs_XM12 vgs_XM12 vds_XM12 cgg_XM12 cgs_XM12 cgd_XM12 cbg_XM12 cbd_XM12 cbs_XM12 cdg_XM12 cdd_XM12 cds_XM12 csg_XM12 csd_XM12 css_XM12 cgb_XM12 cdb_XM12 csb_XM12 cbb_XM12 capbd_XM12 capbs_XM12 gmbs_XM18 gm_XM18 gds_XM18 vdsat_XM18 vth_XM18 id_XM18 ibd_XM18 ibs_XM18 gbd_XM18 gbs_XM18 isub_XM18 igidl_XM18 igisl_XM18 igs_XM18 igd_XM18 igb_XM18 igcs_XM18 vbs_XM18 vgs_XM18 vds_XM18 cgg_XM18 cgs_XM18 cgd_XM18 cbg_XM18 cbd_XM18 cbs_XM18 cdg_XM18 cdd_XM18 cds_XM18 csg_XM18 csd_XM18 css_XM18 cgb_XM18 cdb_XM18 csb_XM18 cbb_XM18 capbd_XM18 capbs_XM18 gmbs_XM13 gm_XM13 gds_XM13 vdsat_XM13 vth_XM13 id_XM13 ibd_XM13 ibs_XM13 gbd_XM13 gbs_XM13 isub_XM13 igidl_XM13 igisl_XM13 igs_XM13 igd_XM13 igb_XM13 igcs_XM13 vbs_XM13 vgs_XM13 vds_XM13 cgg_XM13 cgs_XM13 cgd_XM13 cbg_XM13 cbd_XM13 cbs_XM13 cdg_XM13 cdd_XM13 cds_XM13 csg_XM13 csd_XM13 css_XM13 cgb_XM13 cdb_XM13 csb_XM13 cbb_XM13 capbd_XM13 capbs_XM13 capacitance_XC0 cap_XC0 c_XC0 ic_XC0 temp_XC0 dtemp_XC0 w_XC0 l_XC0 m_XC0 scale_XC0 i_XC0 p_XC0 sens_dc_XC0 sens_real_XC0 sens_imag_XC0 sens_mag_XC0 sens_ph_XC0 sens_cplx_XC0 capacitance_XC1 cap_XC1 c_XC1 ic_XC1 temp_XC1 dtemp_XC1 w_XC1 l_XC1 m_XC1 scale_XC1 i_XC1 p_XC1 sens_dc_XC1 sens_real_XC1 sens_imag_XC1 sens_mag_XC1 sens_ph_XC1 sens_cplx_XC1 
